module and_gate(
	input a,
	input b,
	output c);

and(c,a,b);

endmodule
